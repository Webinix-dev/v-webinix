module vwebinix

#include "@VMODROOT/src/webinix/include/webinix.h"
$if macos {
	#include "@VMODROOT/src/webinix/src/webview/wkwebview.m"
}

#flag -I@VMODROOT/src/webinix/include/ -DNDEBUG -DNO_CACHING -DNO_CGI -DUSE_WEBSOCKET
#flag @VMODROOT/src/webinix/src/civetweb/civetweb.c
#flag @VMODROOT/src/webinix/src/webinix.c

#flag darwin -framework WebKit -framework Cocoa
#flag windows -lWs2_32 -lOle32

$if msvc {
	#flag -lAdvapi32 -lShell32 -lUser32
}
$if use_tls ? {
	#flag -DWEBUI_USE_TLS -DWEBUI_TLS -DNO_SSL_DL -DOPENSSL_API_1_1
	#flag -lssl -lcrypto
	#flag windows -lBcrypt
} $else {
	#flag -DNO_SSL
}
$if webinix_log ? {
	#flag -DWEBUI_LOG
}

@[typedef]
struct C.webinix_event_t {
pub:
	window       Window    // The window object number
	event_type   EventType // Event type
	element      &char     // HTML element ID
	event_number usize     // Internal Webinix
	bind_id      usize     // Bind ID
}

// -- Definitions ---------------------
fn C.webinix_new_window() Window
fn C.webinix_new_window_id(win_id Window)
fn C.webinix_get_new_window_id() Window
fn C.webinix_bind(win Window, elem &char, func fn (&C.webinix_event_t)) Function
fn C.webinix_get_best_browser(win Window) Browser
fn C.webinix_show(win Window, content &char) bool
fn C.webinix_show_browser(win Window, content &char, browser Browser) bool
fn C.webinix_show_wv(win Window, content &char) bool
fn C.webinix_set_kiosk(win Window, kiosk bool)
fn C.webinix_wait()
fn C.webinix_close(win Window)
fn C.webinix_destroy(win Window)
fn C.webinix_exit()
fn C.webinix_set_root_folder(win Window, path &char)
fn C.webinix_set_default_root_folder(path &char)
fn C.webinix_set_file_handler(win Window, handler fn (file_name &char, length int)) // not wrapped
fn C.webinix_is_shown(win Window) bool
fn C.webinix_set_timeout(second usize)
fn C.webinix_set_icon(win Window, icon &char, icon_type &char)
fn C.webinix_encode(str &char) &char
fn C.webinix_decode(str &char) &char
fn C.webinix_free(ptr voidptr) // not wrapped
fn C.webinix_malloc(size usize) voidptr // not wrapped
fn C.webinix_send_raw(size Window, func &char, raw voidptr, size usize) // not wrapped
fn C.webinix_set_hide(win Window, status bool)
fn C.webinix_set_size(win Window, width usize, height usize)
fn C.webinix_set_position(win Window, x usize, y usize)
fn C.webinix_set_profile(win Window, name &char, path &char)
fn C.webinix_set_proxy(win Window, proxy_server &char)
fn C.webinix_get_url(win Window) &char
fn C.webinix_set_public(win Window, status bool)
fn C.webinix_navigate(win Window, url &char)
fn C.webinix_clean()
fn C.webinix_delete_all_profiles()
fn C.webinix_delete_profile(win Window)
fn C.webinix_get_parent_process_id(win Window) usize
fn C.webinix_get_child_process_id(win Window) usize
fn C.webinix_set_port(win Window, port usize) bool
// fn C.webinix_config(option Config, port usize) bool
fn C.webinix_set_tls_certificate(certificate_pem &char, private_key_pem &char) bool

// -- JavaScript ----------------------
fn C.webinix_run(win Window, script &char)
fn C.webinix_script(win Window, script &char, timeout usize, buffer &char, buffer_length usize) bool
fn C.webinix_set_runtime(win Window, runtime Runtime)
fn C.webinix_get_count(e &C.webinix_event_t) usize
fn C.webinix_get_int(e &C.webinix_event_t) i64
fn C.webinix_get_int_at(e &C.webinix_event_t, idx usize) i64
fn C.webinix_get_float(e &C.webinix_event_t) f64
fn C.webinix_get_float_at(e &C.webinix_event_t, idx usize) f64
fn C.webinix_get_string(e &C.webinix_event_t) &char
fn C.webinix_get_string_at(e &C.webinix_event_t, idx usize) &char
fn C.webinix_get_bool(e &C.webinix_event_t) bool
fn C.webinix_get_bool_at(e &C.webinix_event_t, idx usize) bool
fn C.webinix_get_size(e &C.webinix_event_t) usize
fn C.webinix_get_size_at(e &C.webinix_event_t, idx usize) usize
fn C.webinix_return_int(e &C.webinix_event_t, n i64)
fn C.webinix_return_string(e &C.webinix_event_t, s &char)
fn C.webinix_return_bool(e &C.webinix_event_t, b bool)

// -- Interface ----------------------- // not wrapped
fn C.webinix_interface_bind(win Window, element &char, func fn (win Window, event_type EventType, element &char, event_num usize, bind_id usize)) Function
fn C.webinix_interface_set_response(win Window, event_num usize, resp &char)
fn C.webinix_interface_is_app_running() bool
fn C.webinix_interface_get_window_id(win Window) Window
