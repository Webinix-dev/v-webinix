/*
V-Webinix 2.4.0-beta
https://github.com/webinix-dev/v-webinix
Copyright (c) 2023 Mehmet Ali.
Licensed under MIT License.
All rights reserved.
*/

module vwebinix

import json

pub type Window = usize

pub type Function = usize

pub type Event = C.webinix_event_t

[params]
pub struct ScriptOptions {
	max_response_size usize = 8192
	timeout           usize
}

pub enum EventType {
	disconnected        = 0
	connected           = 1
	multi_connection    = 2
	unwanted_connection = 3
	mouse_click         = 4
	navigation          = 5
	callback            = 6
}

pub enum Browser {
	any      = 0
	chrome   = 1
	firefox  = 2
	edge     = 3
	safari   = 4
	chromium = 5
	opera    = 6
	brave    = 7
	vivaldi  = 8
	epic     = 9
	yandex   = 10
}

pub enum Runtime {
	@none  = 0
	deno   = 1
	nodejs = 2
}

// == Definitions =============================================================

// Create a new webinix window object.
pub fn new_window() Window {
	return C.webinix_new_window()
}

// Create a new webinix window object.
pub fn (w Window) new_window() {
	C.webinix_new_window_id(w)
}

// Get a free window ID that can be used with the `new_window` method.
pub fn get_new_window_id() Window {
	return C.webinix_get_new_window_id()
}

// Bind a specific html element click event with a function. Empty element means all events.
pub fn (w Window) bind(element string, func fn (&Event)) Function {
	return C.webinix_bind(w, &char(element.str), func)
}

// Show a window using embedded HTML, or a file. If the window is already open, it will be refreshed.
pub fn (w Window) show(content string) ! {
	if !C.webinix_show(w, &char(content.str)) {
		return error('Failed showing window.')
	}
}

// Show a window using embedded HTML, or a file in a specified browser. If the window is already open, it will be refreshed.
pub fn (w Window) show_browser(content string, browser Browser) ! {
	if !C.webinix_show_browser(w, &char(content.str), browser) {
		return error('Failed showing window in `${browser}`.')
	}
}

// Set the window in Kiosk mode (full screen).
pub fn (w Window) set_kiosk(kiosk bool) {
	C.webinix_set_kiosk(w, kiosk)
}

// Set the web-server root folder path for a specific window.
pub fn (w Window) set_root_folder(path string) {
	C.webinix_set_root_folder(w, &char(path.str))
}

// Set the web-server root folder path for all windows.
pub fn set_root_folder(path string) {
	C.webinix_set_default_root_folder(&char(path.str))
}

// Wait until all opened windows get closed.
pub fn wait() {
	C.webinix_wait()
}

// Close the window. The window object will still exist.
pub fn (w Window) close() {
	C.webinix_close(w)
}

// Close the window and free all memory resources.
pub fn (w Window) destroy() {
	C.webinix_destroy(w)
}

// Close all open windows. `wait()` will break.
pub fn exit() {
	C.webinix_exit()
}

// == Other ===================================================================

// Check if the window is still running.
pub fn (w Window) is_shown() bool {
	return C.webinix_is_shown(w)
}

// Set the maximum time in seconds to wait for the browser to start.
pub fn set_timeout(timeout usize) {
	C.webinix_set_timeout(timeout)
}

// Set the default embedded HTML favicon.
pub fn (w Window) set_icon(icon string, icon_type string) {
	C.webinix_set_icon(w, &char(icon.str), &char(icon_type.str))
}

// Allow the window URL to be re-used in normal web browsers.
pub fn (w Window) set_multi_access(status bool) {
	C.webinix_set_multi_access(w, status)
}

// == Javascript ==============================================================

// Run JavaScript without waiting for the response.
pub fn (w Window) run(script string) {
	C.webinix_run(w, &char(script.str))
}

// Run JavaScript and get the response back (Make sure your local buffer can hold the response).
pub fn (w Window) script(javascript string, opts ScriptOptions) !string {
	mut buffer := []u8{len: int(opts.max_response_size)}.str().str
	if !C.webinix_script(w, &char(javascript.str), opts.timeout, &char(buffer), opts.max_response_size) {
		return error('Failed running script. `${javascript}`')
	}
	return unsafe { buffer.vstring() }
}

// Chose between Deno and Nodejs as runtime for .js and .ts files.
pub fn (w Window) set_runtime(runtime Runtime) {
	C.webinix_set_runtime(w, runtime)
}

// Parse argument as integer.
pub fn (e &Event) int() int {
	return int(C.webinix_get_int(e))
}

// Parse argument as integer.
pub fn (e &Event) i64() i64 {
	return C.webinix_get_int(e)
}

// Parse argument as string.
pub fn (e &Event) string() string {
	// Ensure GCC and Clang compiles with `-cstrict`
	return unsafe { (&char(C.webinix_get_string(e))).vstring() }
}

// Parse argument as boolean.
pub fn (e &Event) bool() bool {
	return C.webinix_get_bool(e)
}

// Decode arguments into a V data type.
pub fn (e Event) decode[T]() !T {
	return json.decode(T, e.string()) or { return error('Failed decoding arguments. `${err}`') }
}

type Response = bool | i64 | int | string

// Return the response to JavaScript.
pub fn (e &Event) @return(response Response) {
	match response {
		int {
			C.webinix_return_int(e, i64(response))
		}
		i64 {
			C.webinix_return_int(e, response)
		}
		string {
			C.webinix_return_string(e, &char(response.str))
		}
		bool {
			C.webinix_return_bool(e, response)
		}
	}
}

// Run the window in hidden mode.
pub fn (w Window) set_hide(status bool) {
	C.webinix_set_hide(w, status)
}

// Set the window size.
pub fn (w Window) set_size(width usize, height usize) {
	C.webinix_set_size(w, width, height)
}

// Set the window position.
pub fn (w Window) set_position(x usize, y usize) {
	C.webinix_set_position(w, x, y)
}
